library ieee;
use ieee.std_logic_1164.all;

entity MIPS is
  port (
    clock : in std_logic;
    reset : in std_logic
  ) ;
end MIPS ;

architecture Behavior of MIPS is

  signal

begin



end architecture ; -- Behavior