library ieee ;
    use ieee.std_logic_1164.all ;
    use ieee.numeric_std.all ;

entity IF_ID is
  port (
    clock
  ) ;
end IF_ID ; 

architecture Behavior of IF_ID is

begin

end architecture ;