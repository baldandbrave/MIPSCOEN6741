library ieee ;
    use ieee.std_logic_1164.all ;
    use ieee.numeric_std.all ;

entity ID_EX is
  port (
    clock
  ) ;
end ID_EX ; 

architecture Behavior of ID_EX is

begin

end architecture ;