library ieee ;
    use ieee.std_logic_1164.all ;
    use ieee.numeric_std.all ;

entity EX_MEM is
  port (
    clock
  ) ;
end EX_MEM ; 

architecture Behavior of EX_MEM is

begin

end architecture ;