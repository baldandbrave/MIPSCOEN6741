library ieee ;
    use ieee.std_logic_1164.all ;
    use ieee.numeric_std.all ;

entity MEM_WB is
  port (
    clock
  ) ;
end MEM_WB ; 

architecture Behavior of MEM_WB is

begin

end architecture ;